`define BUILD_DATE "20230529"
`define XILINX 1
`define LARGE_FPGA 1
`define MISTEX_HDMI 1
`define CLK_100_EXT 1
`define MISTER_DOWNSCALE_NN 1
`define MISTER_DISABLE_YC 1
`define MISTER_DISABLE_ALSA 1
`define SKIP_IIR_FILTER 1
`define MISTER_FB 1
